-------------------------------------------------------------------------------
-- Title : uscite
-- Project :
-------------------------------------------------------------------------------
-- File : uscite.vhd
-- Author : <franc@DESKTOP-5J5ST91>
-- Company :
-- Created : 2020-03-22
-- Last update: 2020-03-22
-- Platform :
-- Standard : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-------------------------------------------------------------------------------
-- Copyright (c) 2020
-------------------------------------------------------------------------------
-- Revisions :
-- Date Version Author Description
-- 2020-03-22 1.0 franc Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity uscite is

port (
OINV : out std_logic;
OAND : out std_logic;
OOR : out std_logic;
OXOR : out std_logic;
IINV : in std_logic;
IAND : in std_logic;
IOR : in std_logic;
IXOR : in std_logic);

end uscite;

-------------------------------------------------------------------------------

architecture str of uscite is

-----------------------------------------------------------------------------
-- Internal signal declarations
-----------------------------------------------------------------------------

begin -- architecture str

OINV <= IINV;
OAND <= IAND;
OOR <= IOR;
OXOR <= IXOR;
-----------------------------------------------------------------------------
-- Component instantiations
-----------------------------------------------------------------------------

end architecture str;

-------------------------------------------------------------------------------
